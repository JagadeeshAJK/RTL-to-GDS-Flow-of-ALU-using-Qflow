module ALU (A[0], A[1], A[2], A[3], A[4], A[5], A[6], A[7], B[0], B[1], B[2], B[3], B[4], B[5], B[6], B[7], select[0], select[1], select[2], select[3], clk, ALU_out[0], ALU_out[1], ALU_out[2], ALU_out[3], ALU_out[4], ALU_out[5], ALU_out[6], ALU_out[7], Carry_out);

input A[0];
input A[1];
input A[2];
input A[3];
input A[4];
input A[5];
input A[6];
input A[7];
input B[0];
input B[1];
input B[2];
input B[3];
input B[4];
input B[5];
input B[6];
input B[7];
input select[0];
input select[1];
input select[2];
input select[3];
input clk;
output ALU_out[0];
output ALU_out[1];
output ALU_out[2];
output ALU_out[3];
output ALU_out[4];
output ALU_out[5];
output ALU_out[6];
output ALU_out[7];
output Carry_out;

BUFX2 BUFX2_1 ( .A(B[1]), .Y(B_1_bF_buf3_) );
BUFX2 BUFX2_2 ( .A(B[1]), .Y(B_1_bF_buf2_) );
BUFX2 BUFX2_3 ( .A(B[1]), .Y(B_1_bF_buf1_) );
BUFX2 BUFX2_4 ( .A(B[1]), .Y(B_1_bF_buf0_) );
BUFX2 BUFX2_5 ( .A(_299_), .Y(_299__bF_buf3) );
BUFX2 BUFX2_6 ( .A(_299_), .Y(_299__bF_buf2) );
BUFX2 BUFX2_7 ( .A(_299_), .Y(_299__bF_buf1) );
BUFX2 BUFX2_8 ( .A(_299_), .Y(_299__bF_buf0) );
BUFX2 BUFX2_9 ( .A(_387_), .Y(_387__bF_buf3) );
BUFX2 BUFX2_10 ( .A(_387_), .Y(_387__bF_buf2) );
BUFX2 BUFX2_11 ( .A(_387_), .Y(_387__bF_buf1) );
BUFX2 BUFX2_12 ( .A(_387_), .Y(_387__bF_buf0) );
BUFX2 BUFX2_13 ( .A(_486_), .Y(_486__bF_buf3) );
BUFX2 BUFX2_14 ( .A(_486_), .Y(_486__bF_buf2) );
BUFX2 BUFX2_15 ( .A(_486_), .Y(_486__bF_buf1) );
BUFX2 BUFX2_16 ( .A(_486_), .Y(_486__bF_buf0) );
BUFX2 BUFX2_17 ( .A(B[2]), .Y(B_2_bF_buf3_) );
BUFX4 BUFX4_1 ( .A(B[2]), .Y(B_2_bF_buf2_) );
BUFX2 BUFX2_18 ( .A(B[2]), .Y(B_2_bF_buf1_) );
BUFX2 BUFX2_19 ( .A(B[2]), .Y(B_2_bF_buf0_) );
NAND2X1 NAND2X1_1 ( .A(_105_), .B(_107_), .Y(_108_) );
NAND3X1 NAND3X1_1 ( .A(_354_), .B(_108_), .C(_103_), .Y(_109_) );
OAI21X1 OAI21X1_1 ( .A(A[3]), .B(_92_), .C(_109_), .Y(_110_) );
OAI21X1 OAI21X1_2 ( .A(_812_), .B(_45_), .C(_657_), .Y(_111_) );
INVX1 INVX1_1 ( .A(_111_), .Y(_112_) );
AOI21X1 AOI21X1_1 ( .A(_103_), .B(_354_), .C(_112_), .Y(_113_) );
OAI21X1 OAI21X1_3 ( .A(_668_), .B(_113_), .C(_409_), .Y(_114_) );
NAND2X1 NAND2X1_2 ( .A(_67_), .B(_68_), .Y(_115_) );
NAND2X1 NAND2X1_3 ( .A(B[0]), .B(_679_), .Y(_116_) );
OAI21X1 OAI21X1_4 ( .A(_116_), .B(_56_), .C(A[4]), .Y(_117_) );
INVX1 INVX1_2 ( .A(_116_), .Y(_118_) );
NAND3X1 NAND3X1_2 ( .A(_79_), .B(_118_), .C(_28_), .Y(_119_) );
AOI21X1 AOI21X1_2 ( .A(_117_), .B(_119_), .C(B_1_bF_buf3_), .Y(_120_) );
AOI21X1 AOI21X1_3 ( .A(_86_), .B(_88_), .C(_120_), .Y(_121_) );
OAI21X1 OAI21X1_5 ( .A(_76_), .B(_121_), .C(_78_), .Y(_122_) );
NAND2X1 NAND2X1_4 ( .A(_115_), .B(_122_), .Y(_123_) );
INVX1 INVX1_3 ( .A(_115_), .Y(_124_) );
INVX1 INVX1_4 ( .A(_93_), .Y(_125_) );
NAND3X1 NAND3X1_3 ( .A(_86_), .B(_101_), .C(_95_), .Y(_126_) );
NAND3X1 NAND3X1_4 ( .A(_124_), .B(_125_), .C(_126_), .Y(_127_) );
NAND2X1 NAND2X1_5 ( .A(_127_), .B(_123_), .Y(_128_) );
NAND2X1 NAND2X1_6 ( .A(_92_), .B(_128_), .Y(_129_) );
OAI21X1 OAI21X1_6 ( .A(_51_), .B(_45_), .C(_49_), .Y(_130_) );
AOI21X1 AOI21X1_4 ( .A(_122_), .B(_69_), .C(_59_), .Y(_131_) );
OAI21X1 OAI21X1_7 ( .A(_365_), .B(_131_), .C(_130_), .Y(_132_) );
NAND3X1 NAND3X1_5 ( .A(_376_), .B(_132_), .C(_129_), .Y(_133_) );
OAI21X1 OAI21X1_8 ( .A(_365_), .B(_131_), .C(_111_), .Y(_134_) );
NAND3X1 NAND3X1_6 ( .A(B[5]), .B(_657_), .C(_134_), .Y(_135_) );
NAND2X1 NAND2X1_7 ( .A(_114_), .B(_135_), .Y(_136_) );
OAI21X1 OAI21X1_9 ( .A(_133_), .B(_136_), .C(_114_), .Y(_137_) );
NAND3X1 NAND3X1_7 ( .A(_123_), .B(_127_), .C(_92_), .Y(_138_) );
INVX1 INVX1_5 ( .A(_130_), .Y(_139_) );
OAI21X1 OAI21X1_10 ( .A(_365_), .B(_131_), .C(_139_), .Y(_140_) );
NAND3X1 NAND3X1_8 ( .A(B[4]), .B(_140_), .C(_138_), .Y(_141_) );
NAND2X1 NAND2X1_8 ( .A(_133_), .B(_141_), .Y(_142_) );
NOR2X1 NOR2X1_1 ( .A(_136_), .B(_142_), .Y(_143_) );
OAI21X1 OAI21X1_11 ( .A(_74_), .B(_45_), .C(_98_), .Y(_144_) );
INVX1 INVX1_6 ( .A(_144_), .Y(_145_) );
OAI21X1 OAI21X1_12 ( .A(_365_), .B(_131_), .C(_145_), .Y(_146_) );
XOR2X1 XOR2X1_1 ( .A(_121_), .B(_101_), .Y(_147_) );
NAND2X1 NAND2X1_9 ( .A(_147_), .B(_92_), .Y(_148_) );
NAND3X1 NAND3X1_9 ( .A(_431_), .B(_146_), .C(_148_), .Y(_149_) );
XOR2X1 XOR2X1_2 ( .A(_95_), .B(_85_), .Y(_150_) );
NAND3X1 NAND3X1_10 ( .A(_354_), .B(_150_), .C(_103_), .Y(_151_) );
OAI21X1 OAI21X1_13 ( .A(_365_), .B(_131_), .C(_87_), .Y(_152_) );
NAND3X1 NAND3X1_11 ( .A(_486__bF_buf3), .B(_151_), .C(_152_), .Y(_153_) );
OAI21X1 OAI21X1_14 ( .A(_365_), .B(_131_), .C(_144_), .Y(_154_) );
INVX1 INVX1_7 ( .A(_147_), .Y(_155_) );
NAND2X1 NAND2X1_10 ( .A(_155_), .B(_92_), .Y(_156_) );
NAND3X1 NAND3X1_12 ( .A(B[3]), .B(_154_), .C(_156_), .Y(_157_) );
NAND2X1 NAND2X1_11 ( .A(_149_), .B(_157_), .Y(_158_) );
OAI21X1 OAI21X1_15 ( .A(_153_), .B(_158_), .C(_149_), .Y(_159_) );
AOI21X1 AOI21X1_5 ( .A(_143_), .B(_159_), .C(_137_), .Y(_160_) );
OAI21X1 OAI21X1_16 ( .A(_365_), .B(_131_), .C(_104_), .Y(_161_) );
NAND3X1 NAND3X1_13 ( .A(_387__bF_buf3), .B(_109_), .C(_161_), .Y(_162_) );
AOI21X1 AOI21X1_6 ( .A(_161_), .B(_109_), .C(_387__bF_buf2), .Y(_163_) );
NOR2X1 NOR2X1_2 ( .A(A[2]), .B(_299__bF_buf3), .Y(_164_) );
OAI21X1 OAI21X1_17 ( .A(_164_), .B(_163_), .C(_162_), .Y(_165_) );
INVX1 INVX1_8 ( .A(_87_), .Y(_166_) );
OAI21X1 OAI21X1_18 ( .A(_365_), .B(_131_), .C(_166_), .Y(_167_) );
XOR2X1 XOR2X1_3 ( .A(_95_), .B(_86_), .Y(_168_) );
NAND3X1 NAND3X1_14 ( .A(_354_), .B(_168_), .C(_103_), .Y(_169_) );
NAND3X1 NAND3X1_15 ( .A(B_2_bF_buf3_), .B(_169_), .C(_167_), .Y(_170_) );
NAND2X1 NAND2X1_12 ( .A(_153_), .B(_170_), .Y(_171_) );
NOR2X1 NOR2X1_3 ( .A(_171_), .B(_158_), .Y(_172_) );
NAND3X1 NAND3X1_16 ( .A(_165_), .B(_172_), .C(_143_), .Y(_173_) );
AOI21X1 AOI21X1_7 ( .A(_160_), .B(_173_), .C(_343_), .Y(_174_) );
NAND2X1 NAND2X1_13 ( .A(B_1_bF_buf2_), .B(_110_), .Y(_175_) );
NAND2X1 NAND2X1_14 ( .A(_162_), .B(_175_), .Y(_176_) );
XOR2X1 XOR2X1_4 ( .A(_176_), .B(_164_), .Y(_177_) );
NAND2X1 NAND2X1_15 ( .A(_177_), .B(_174_), .Y(_178_) );
OAI21X1 OAI21X1_19 ( .A(_110_), .B(_174_), .C(_178_), .Y(_179_) );
NAND3X1 NAND3X1_17 ( .A(B[0]), .B(_354_), .C(_103_), .Y(_180_) );
NAND2X1 NAND2X1_16 ( .A(A[3]), .B(_180_), .Y(_181_) );
NAND2X1 NAND2X1_17 ( .A(_85_), .B(_92_), .Y(_182_) );
AOI21X1 AOI21X1_8 ( .A(_181_), .B(_182_), .C(B_1_bF_buf1_), .Y(_183_) );
INVX1 INVX1_9 ( .A(_164_), .Y(_184_) );
AOI21X1 AOI21X1_9 ( .A(_175_), .B(_184_), .C(_183_), .Y(_185_) );
OAI21X1 OAI21X1_20 ( .A(_171_), .B(_185_), .C(_153_), .Y(_186_) );
AND2X2 AND2X2_1 ( .A(_149_), .B(_157_), .Y(_187_) );
NOR2X1 NOR2X1_4 ( .A(_187_), .B(_186_), .Y(_188_) );
AND2X2 AND2X2_2 ( .A(_186_), .B(_187_), .Y(_189_) );
OAI21X1 OAI21X1_21 ( .A(_188_), .B(_189_), .C(_174_), .Y(_190_) );
OAI21X1 OAI21X1_22 ( .A(_144_), .B(_92_), .C(_148_), .Y(_191_) );
INVX1 INVX1_10 ( .A(_149_), .Y(_192_) );
INVX1 INVX1_11 ( .A(_153_), .Y(_193_) );
AOI21X1 AOI21X1_10 ( .A(_193_), .B(_157_), .C(_192_), .Y(_194_) );
NAND3X1 NAND3X1_18 ( .A(_486__bF_buf2), .B(_169_), .C(_167_), .Y(_195_) );
NAND3X1 NAND3X1_19 ( .A(B_2_bF_buf2_), .B(_151_), .C(_152_), .Y(_196_) );
NAND2X1 NAND2X1_18 ( .A(_195_), .B(_196_), .Y(_197_) );
NAND3X1 NAND3X1_20 ( .A(_149_), .B(_157_), .C(_197_), .Y(_198_) );
OAI21X1 OAI21X1_23 ( .A(_185_), .B(_198_), .C(_194_), .Y(_199_) );
AOI21X1 AOI21X1_11 ( .A(_199_), .B(_143_), .C(_137_), .Y(_200_) );
OAI21X1 OAI21X1_24 ( .A(_343_), .B(_200_), .C(_191_), .Y(_201_) );
AOI21X1 AOI21X1_12 ( .A(_190_), .B(_201_), .C(_376_), .Y(_202_) );
INVX1 INVX1_12 ( .A(_137_), .Y(_203_) );
NAND2X1 NAND2X1_19 ( .A(_159_), .B(_143_), .Y(_204_) );
NAND3X1 NAND3X1_21 ( .A(_203_), .B(_204_), .C(_173_), .Y(_205_) );
XOR2X1 XOR2X1_5 ( .A(_165_), .B(_197_), .Y(_206_) );
INVX1 INVX1_13 ( .A(_206_), .Y(_207_) );
NAND3X1 NAND3X1_22 ( .A(_332_), .B(_207_), .C(_205_), .Y(_208_) );
OAI21X1 OAI21X1_25 ( .A(_166_), .B(_92_), .C(_151_), .Y(_209_) );
OAI21X1 OAI21X1_26 ( .A(_343_), .B(_200_), .C(_209_), .Y(_210_) );
NAND3X1 NAND3X1_23 ( .A(_431_), .B(_208_), .C(_210_), .Y(_212_) );
NAND3X1 NAND3X1_24 ( .A(_376_), .B(_201_), .C(_190_), .Y(_213_) );
OAI21X1 OAI21X1_27 ( .A(_212_), .B(_202_), .C(_213_), .Y(_214_) );
NAND3X1 NAND3X1_25 ( .A(_197_), .B(_187_), .C(_165_), .Y(_215_) );
AOI21X1 AOI21X1_13 ( .A(_215_), .B(_194_), .C(_142_), .Y(_216_) );
NAND3X1 NAND3X1_26 ( .A(_142_), .B(_194_), .C(_215_), .Y(_217_) );
INVX1 INVX1_14 ( .A(_217_), .Y(_218_) );
OAI21X1 OAI21X1_28 ( .A(_216_), .B(_218_), .C(_174_), .Y(_219_) );
OAI21X1 OAI21X1_29 ( .A(_139_), .B(_92_), .C(_129_), .Y(_220_) );
OAI21X1 OAI21X1_30 ( .A(_343_), .B(_200_), .C(_220_), .Y(_221_) );
NAND3X1 NAND3X1_27 ( .A(_409_), .B(_221_), .C(_219_), .Y(_223_) );
OAI21X1 OAI21X1_31 ( .A(_112_), .B(_92_), .C(_657_), .Y(_224_) );
INVX1 INVX1_15 ( .A(_224_), .Y(_225_) );
AOI21X1 AOI21X1_14 ( .A(_205_), .B(_332_), .C(_225_), .Y(_226_) );
OAI21X1 OAI21X1_32 ( .A(_668_), .B(_226_), .C(_398_), .Y(_227_) );
OAI21X1 OAI21X1_33 ( .A(_343_), .B(_200_), .C(_224_), .Y(_228_) );
NAND3X1 NAND3X1_28 ( .A(B[6]), .B(_657_), .C(_228_), .Y(_229_) );
NAND2X1 NAND2X1_20 ( .A(_229_), .B(_227_), .Y(_230_) );
OAI21X1 OAI21X1_34 ( .A(_223_), .B(_230_), .C(_227_), .Y(_231_) );
INVX1 INVX1_16 ( .A(_216_), .Y(_232_) );
NAND3X1 NAND3X1_29 ( .A(_232_), .B(_217_), .C(_174_), .Y(_234_) );
INVX1 INVX1_17 ( .A(_220_), .Y(_235_) );
OAI21X1 OAI21X1_35 ( .A(_343_), .B(_200_), .C(_235_), .Y(_236_) );
NAND3X1 NAND3X1_30 ( .A(B[5]), .B(_236_), .C(_234_), .Y(_237_) );
NAND2X1 NAND2X1_21 ( .A(_223_), .B(_237_), .Y(_238_) );
NOR2X1 NOR2X1_5 ( .A(_230_), .B(_238_), .Y(_239_) );
AOI21X1 AOI21X1_15 ( .A(_239_), .B(_214_), .C(_231_), .Y(_240_) );
INVX1 INVX1_18 ( .A(_110_), .Y(_241_) );
OAI21X1 OAI21X1_36 ( .A(_343_), .B(_200_), .C(_241_), .Y(_242_) );
AOI21X1 AOI21X1_16 ( .A(_178_), .B(_242_), .C(B_2_bF_buf1_), .Y(_243_) );
INVX1 INVX1_19 ( .A(_243_), .Y(_245_) );
NAND3X1 NAND3X1_31 ( .A(B_2_bF_buf0_), .B(_242_), .C(_178_), .Y(_246_) );
INVX2 INVX2_1 ( .A(A[2]), .Y(_247_) );
NOR2X1 NOR2X1_6 ( .A(B[0]), .B(_247_), .Y(_248_) );
NOR2X1 NOR2X1_7 ( .A(_164_), .B(_248_), .Y(_249_) );
NAND3X1 NAND3X1_32 ( .A(_332_), .B(_249_), .C(_205_), .Y(_250_) );
OAI21X1 OAI21X1_37 ( .A(_343_), .B(_200_), .C(_247_), .Y(_251_) );
NAND3X1 NAND3X1_33 ( .A(_387__bF_buf1), .B(_250_), .C(_251_), .Y(_252_) );
NOR2X1 NOR2X1_8 ( .A(A[1]), .B(_299__bF_buf2), .Y(_253_) );
AOI21X1 AOI21X1_17 ( .A(_251_), .B(_250_), .C(_387__bF_buf0), .Y(_254_) );
OAI21X1 OAI21X1_38 ( .A(_253_), .B(_254_), .C(_252_), .Y(_256_) );
NAND2X1 NAND2X1_22 ( .A(_246_), .B(_256_), .Y(_257_) );
NAND2X1 NAND2X1_23 ( .A(_245_), .B(_257_), .Y(_258_) );
NAND3X1 NAND3X1_34 ( .A(_332_), .B(_206_), .C(_205_), .Y(_259_) );
INVX1 INVX1_20 ( .A(_209_), .Y(_260_) );
OAI21X1 OAI21X1_39 ( .A(_343_), .B(_200_), .C(_260_), .Y(_261_) );
NAND3X1 NAND3X1_35 ( .A(B[3]), .B(_259_), .C(_261_), .Y(_262_) );
NAND2X1 NAND2X1_24 ( .A(_212_), .B(_262_), .Y(_263_) );
NAND2X1 NAND2X1_25 ( .A(_201_), .B(_190_), .Y(_264_) );
NAND2X1 NAND2X1_26 ( .A(B[4]), .B(_264_), .Y(_265_) );
NAND2X1 NAND2X1_27 ( .A(_213_), .B(_265_), .Y(_267_) );
NOR2X1 NOR2X1_9 ( .A(_263_), .B(_267_), .Y(_268_) );
NAND3X1 NAND3X1_36 ( .A(_268_), .B(_239_), .C(_258_), .Y(_269_) );
AOI21X1 AOI21X1_18 ( .A(_269_), .B(_240_), .C(B[7]), .Y(_270_) );
AOI21X1 AOI21X1_19 ( .A(_256_), .B(_246_), .C(_243_), .Y(_271_) );
AND2X2 AND2X2_3 ( .A(_212_), .B(_262_), .Y(_272_) );
INVX1 INVX1_21 ( .A(_213_), .Y(_273_) );
NOR2X1 NOR2X1_10 ( .A(_202_), .B(_273_), .Y(_274_) );
NAND3X1 NAND3X1_37 ( .A(_272_), .B(_274_), .C(_239_), .Y(_275_) );
OAI21X1 OAI21X1_40 ( .A(_271_), .B(_275_), .C(_240_), .Y(_276_) );
NAND2X1 NAND2X1_28 ( .A(_246_), .B(_245_), .Y(_278_) );
XOR2X1 XOR2X1_6 ( .A(_278_), .B(_256_), .Y(_279_) );
NAND3X1 NAND3X1_38 ( .A(_464_), .B(_279_), .C(_276_), .Y(_280_) );
OAI21X1 OAI21X1_41 ( .A(_179_), .B(_270_), .C(_280_), .Y(_281_) );
OAI21X1 OAI21X1_42 ( .A(B[3]), .B(_281_), .C(_321_), .Y(_282_) );
NAND2X1 NAND2X1_29 ( .A(B[3]), .B(_281_), .Y(_283_) );
OAI21X1 OAI21X1_43 ( .A(A[2]), .B(_174_), .C(_250_), .Y(_284_) );
INVX1 INVX1_22 ( .A(_284_), .Y(_285_) );
INVX1 INVX1_23 ( .A(_253_), .Y(_286_) );
NAND2X1 NAND2X1_30 ( .A(B_1_bF_buf0_), .B(_284_), .Y(_287_) );
NAND3X1 NAND3X1_39 ( .A(_252_), .B(_286_), .C(_287_), .Y(_289_) );
INVX1 INVX1_24 ( .A(_252_), .Y(_290_) );
OAI21X1 OAI21X1_44 ( .A(_254_), .B(_290_), .C(_253_), .Y(_291_) );
NAND2X1 NAND2X1_31 ( .A(_289_), .B(_291_), .Y(_292_) );
NAND3X1 NAND3X1_40 ( .A(_464_), .B(_292_), .C(_276_), .Y(_293_) );
OAI21X1 OAI21X1_45 ( .A(_285_), .B(_270_), .C(_293_), .Y(_294_) );
NAND2X1 NAND2X1_32 ( .A(B_2_bF_buf3_), .B(_294_), .Y(_295_) );
INVX1 INVX1_25 ( .A(_292_), .Y(_296_) );
NAND3X1 NAND3X1_41 ( .A(_464_), .B(_296_), .C(_276_), .Y(_297_) );
OAI21X1 OAI21X1_46 ( .A(_284_), .B(_270_), .C(_297_), .Y(_298_) );
NAND2X1 NAND2X1_33 ( .A(_464_), .B(_276_), .Y(_300_) );
OAI21X1 OAI21X1_47 ( .A(_299__bF_buf1), .B(_300_), .C(A[1]), .Y(_301_) );
NOR2X1 NOR2X1_11 ( .A(B_1_bF_buf3_), .B(_310_), .Y(_302_) );
AOI21X1 AOI21X1_20 ( .A(_270_), .B(_253_), .C(_302_), .Y(_303_) );
AOI22X1 AOI22X1_1 ( .A(_298_), .B(_486__bF_buf1), .C(_301_), .D(_303_), .Y(_304_) );
NAND3X1 NAND3X1_42 ( .A(_283_), .B(_295_), .C(_304_), .Y(_305_) );
INVX1 INVX1_26 ( .A(_179_), .Y(_306_) );
INVX1 INVX1_27 ( .A(_212_), .Y(_307_) );
AOI21X1 AOI21X1_21 ( .A(_265_), .B(_307_), .C(_273_), .Y(_308_) );
INVX1 INVX1_28 ( .A(_223_), .Y(_309_) );
INVX1 INVX1_29 ( .A(_227_), .Y(_311_) );
AOI21X1 AOI21X1_22 ( .A(_309_), .B(_229_), .C(_311_), .Y(_312_) );
AND2X2 AND2X2_4 ( .A(_237_), .B(_223_), .Y(_313_) );
AND2X2 AND2X2_5 ( .A(_227_), .B(_229_), .Y(_314_) );
NAND2X1 NAND2X1_34 ( .A(_314_), .B(_313_), .Y(_315_) );
OAI21X1 OAI21X1_48 ( .A(_308_), .B(_315_), .C(_312_), .Y(_316_) );
NAND3X1 NAND3X1_43 ( .A(_213_), .B(_265_), .C(_272_), .Y(_317_) );
NOR2X1 NOR2X1_12 ( .A(_317_), .B(_315_), .Y(_318_) );
AOI21X1 AOI21X1_23 ( .A(_318_), .B(_258_), .C(_316_), .Y(_319_) );
OAI21X1 OAI21X1_49 ( .A(B[7]), .B(_319_), .C(_306_), .Y(_320_) );
NAND3X1 NAND3X1_44 ( .A(_431_), .B(_280_), .C(_320_), .Y(_322_) );
INVX1 INVX1_30 ( .A(_322_), .Y(_323_) );
NOR2X1 NOR2X1_13 ( .A(B_2_bF_buf2_), .B(_294_), .Y(_324_) );
AOI21X1 AOI21X1_24 ( .A(_324_), .B(_283_), .C(_323_), .Y(_325_) );
OAI21X1 OAI21X1_50 ( .A(_282_), .B(_305_), .C(_325_), .Y(_326_) );
OAI21X1 OAI21X1_51 ( .A(_225_), .B(_174_), .C(_657_), .Y(_327_) );
AOI21X1 AOI21X1_25 ( .A(_300_), .B(_327_), .C(_668_), .Y(_328_) );
NOR2X1 NOR2X1_14 ( .A(B[7]), .B(_328_), .Y(_329_) );
NAND3X1 NAND3X1_45 ( .A(_219_), .B(_221_), .C(_300_), .Y(_330_) );
OAI21X1 OAI21X1_52 ( .A(_317_), .B(_271_), .C(_308_), .Y(_331_) );
NAND2X1 NAND2X1_35 ( .A(_313_), .B(_331_), .Y(_333_) );
NAND2X1 NAND2X1_36 ( .A(_268_), .B(_258_), .Y(_334_) );
NAND3X1 NAND3X1_46 ( .A(_238_), .B(_308_), .C(_334_), .Y(_335_) );
NAND3X1 NAND3X1_47 ( .A(_333_), .B(_335_), .C(_270_), .Y(_336_) );
AOI21X1 AOI21X1_26 ( .A(_330_), .B(_336_), .C(B[6]), .Y(_337_) );
OAI21X1 OAI21X1_53 ( .A(_668_), .B(_226_), .C(B[7]), .Y(_338_) );
OAI21X1 OAI21X1_54 ( .A(B[7]), .B(_319_), .C(_327_), .Y(_339_) );
NAND3X1 NAND3X1_48 ( .A(_464_), .B(_657_), .C(_339_), .Y(_340_) );
NAND2X1 NAND2X1_37 ( .A(_338_), .B(_340_), .Y(_341_) );
AOI21X1 AOI21X1_27 ( .A(_341_), .B(_337_), .C(_329_), .Y(_342_) );
NAND2X1 NAND2X1_38 ( .A(_333_), .B(_335_), .Y(_344_) );
NAND2X1 NAND2X1_39 ( .A(_270_), .B(_344_), .Y(_345_) );
NAND3X1 NAND3X1_49 ( .A(_234_), .B(_236_), .C(_300_), .Y(_346_) );
NAND3X1 NAND3X1_50 ( .A(_398_), .B(_346_), .C(_345_), .Y(_347_) );
NAND3X1 NAND3X1_51 ( .A(B[6]), .B(_336_), .C(_330_), .Y(_348_) );
NAND3X1 NAND3X1_52 ( .A(_348_), .B(_347_), .C(_341_), .Y(_349_) );
INVX1 INVX1_31 ( .A(_264_), .Y(_350_) );
OAI21X1 OAI21X1_55 ( .A(B[7]), .B(_319_), .C(_350_), .Y(_351_) );
OAI21X1 OAI21X1_56 ( .A(_263_), .B(_271_), .C(_212_), .Y(_352_) );
NOR2X1 NOR2X1_15 ( .A(_267_), .B(_352_), .Y(_353_) );
NAND3X1 NAND3X1_53 ( .A(_245_), .B(_252_), .C(_289_), .Y(_355_) );
NAND3X1 NAND3X1_54 ( .A(_246_), .B(_272_), .C(_355_), .Y(_356_) );
AOI21X1 AOI21X1_28 ( .A(_356_), .B(_212_), .C(_274_), .Y(_357_) );
OAI21X1 OAI21X1_57 ( .A(_353_), .B(_357_), .C(_270_), .Y(_358_) );
AOI21X1 AOI21X1_29 ( .A(_358_), .B(_351_), .C(B[5]), .Y(_359_) );
NAND3X1 NAND3X1_55 ( .A(B[5]), .B(_351_), .C(_358_), .Y(_360_) );
OAI21X1 OAI21X1_58 ( .A(_260_), .B(_174_), .C(_208_), .Y(_361_) );
INVX1 INVX1_32 ( .A(_361_), .Y(_362_) );
OAI21X1 OAI21X1_59 ( .A(B[7]), .B(_319_), .C(_362_), .Y(_363_) );
NAND2X1 NAND2X1_40 ( .A(_263_), .B(_271_), .Y(_364_) );
NAND2X1 NAND2X1_41 ( .A(_356_), .B(_364_), .Y(_366_) );
INVX1 INVX1_33 ( .A(_366_), .Y(_367_) );
NAND2X1 NAND2X1_42 ( .A(_367_), .B(_270_), .Y(_368_) );
AOI21X1 AOI21X1_30 ( .A(_368_), .B(_363_), .C(B[4]), .Y(_369_) );
AOI21X1 AOI21X1_31 ( .A(_360_), .B(_369_), .C(_359_), .Y(_370_) );
OAI21X1 OAI21X1_60 ( .A(_370_), .B(_349_), .C(_342_), .Y(_371_) );
OAI21X1 OAI21X1_61 ( .A(B[7]), .B(_319_), .C(_264_), .Y(_372_) );
AOI21X1 AOI21X1_32 ( .A(_356_), .B(_212_), .C(_267_), .Y(_373_) );
NOR2X1 NOR2X1_16 ( .A(_274_), .B(_352_), .Y(_374_) );
OAI21X1 OAI21X1_62 ( .A(_373_), .B(_374_), .C(_270_), .Y(_375_) );
AOI21X1 AOI21X1_33 ( .A(_375_), .B(_372_), .C(B[5]), .Y(_377_) );
AOI21X1 AOI21X1_34 ( .A(_358_), .B(_351_), .C(_409_), .Y(_378_) );
NAND2X1 NAND2X1_43 ( .A(_366_), .B(_270_), .Y(_379_) );
OAI21X1 OAI21X1_63 ( .A(B[7]), .B(_319_), .C(_361_), .Y(_380_) );
AOI21X1 AOI21X1_35 ( .A(_379_), .B(_380_), .C(B[4]), .Y(_381_) );
AOI21X1 AOI21X1_36 ( .A(_368_), .B(_363_), .C(_376_), .Y(_382_) );
OAI22X1 OAI22X1_1 ( .A(_381_), .B(_382_), .C(_377_), .D(_378_), .Y(_383_) );
NOR2X1 NOR2X1_17 ( .A(_383_), .B(_349_), .Y(_384_) );
AOI21X1 AOI21X1_37 ( .A(_384_), .B(_326_), .C(_371_), .Y(_385_) );
OAI21X1 OAI21X1_64 ( .A(B[7]), .B(A[7]), .C(_338_), .Y(_386_) );
INVX1 INVX1_34 ( .A(_386_), .Y(_388_) );
INVX2 INVX2_2 ( .A(A[6]), .Y(_389_) );
NOR2X1 NOR2X1_18 ( .A(B[6]), .B(_389_), .Y(_390_) );
AOI22X1 AOI22X1_2 ( .A(_464_), .B(A[7]), .C(_386_), .D(_390_), .Y(_391_) );
NOR2X1 NOR2X1_19 ( .A(_398_), .B(_389_), .Y(_392_) );
NOR2X1 NOR2X1_20 ( .A(B[6]), .B(A[6]), .Y(_393_) );
INVX2 INVX2_3 ( .A(A[1]), .Y(_394_) );
NOR2X1 NOR2X1_21 ( .A(_387__bF_buf3), .B(_394_), .Y(_395_) );
NOR2X1 NOR2X1_22 ( .A(B_1_bF_buf2_), .B(A[1]), .Y(_396_) );
NOR2X1 NOR2X1_23 ( .A(_396_), .B(_395_), .Y(_397_) );
INVX1 INVX1_35 ( .A(_397_), .Y(_399_) );
OAI21X1 OAI21X1_65 ( .A(_299__bF_buf0), .B(A[0]), .C(_399_), .Y(_400_) );
OAI21X1 OAI21X1_66 ( .A(B_1_bF_buf1_), .B(_394_), .C(_400_), .Y(_401_) );
NOR2X1 NOR2X1_24 ( .A(_486__bF_buf0), .B(_247_), .Y(_402_) );
NOR2X1 NOR2X1_25 ( .A(B_2_bF_buf1_), .B(A[2]), .Y(_403_) );
OAI21X1 OAI21X1_67 ( .A(_402_), .B(_403_), .C(_401_), .Y(_404_) );
OAI21X1 OAI21X1_68 ( .A(B_2_bF_buf0_), .B(_247_), .C(_404_), .Y(_405_) );
OAI21X1 OAI21X1_69 ( .A(_431_), .B(A[3]), .C(_405_), .Y(_406_) );
OAI21X1 OAI21X1_70 ( .A(B[3]), .B(_104_), .C(_406_), .Y(_407_) );
NOR2X1 NOR2X1_26 ( .A(_376_), .B(_79_), .Y(_408_) );
NOR2X1 NOR2X1_27 ( .A(B[4]), .B(A[4]), .Y(_410_) );
OAI21X1 OAI21X1_71 ( .A(_408_), .B(_410_), .C(_407_), .Y(_411_) );
OAI21X1 OAI21X1_72 ( .A(B[4]), .B(_79_), .C(_411_), .Y(_412_) );
OAI21X1 OAI21X1_73 ( .A(_409_), .B(A[5]), .C(_412_), .Y(_413_) );
OAI21X1 OAI21X1_74 ( .A(B[5]), .B(_21_), .C(_413_), .Y(_414_) );
OAI21X1 OAI21X1_75 ( .A(_392_), .B(_393_), .C(_414_), .Y(_415_) );
OAI21X1 OAI21X1_76 ( .A(_415_), .B(_388_), .C(_391_), .Y(_416_) );
NOR2X1 NOR2X1_28 ( .A(select[0]), .B(_233_), .Y(_417_) );
INVX1 INVX1_36 ( .A(select[3]), .Y(_418_) );
INVX1 INVX1_37 ( .A(select[2]), .Y(_419_) );
NOR2X1 NOR2X1_29 ( .A(_418_), .B(_419_), .Y(_421_) );
NAND2X1 NAND2X1_44 ( .A(_417_), .B(_421_), .Y(_422_) );
NOR2X1 NOR2X1_30 ( .A(_431_), .B(_104_), .Y(_423_) );
NOR2X1 NOR2X1_31 ( .A(B[3]), .B(A[3]), .Y(_424_) );
NOR2X1 NOR2X1_32 ( .A(_424_), .B(_423_), .Y(_425_) );
INVX1 INVX1_38 ( .A(_425_), .Y(_426_) );
INVX2 INVX2_4 ( .A(A[0]), .Y(_427_) );
NOR2X1 NOR2X1_33 ( .A(_299__bF_buf3), .B(_427_), .Y(_428_) );
NOR2X1 NOR2X1_34 ( .A(B[0]), .B(A[0]), .Y(_429_) );
NOR2X1 NOR2X1_35 ( .A(_429_), .B(_428_), .Y(_430_) );
INVX1 INVX1_39 ( .A(_430_), .Y(_432_) );
NAND3X1 NAND3X1_56 ( .A(_399_), .B(_426_), .C(_432_), .Y(_433_) );
NOR2X1 NOR2X1_36 ( .A(_393_), .B(_392_), .Y(_434_) );
INVX1 INVX1_40 ( .A(_434_), .Y(_435_) );
NOR2X1 NOR2X1_37 ( .A(_410_), .B(_408_), .Y(_436_) );
INVX2 INVX2_5 ( .A(_436_), .Y(_437_) );
NOR2X1 NOR2X1_38 ( .A(_403_), .B(_402_), .Y(_438_) );
NOR2X1 NOR2X1_39 ( .A(_409_), .B(_21_), .Y(_439_) );
NOR2X1 NOR2X1_40 ( .A(B[5]), .B(A[5]), .Y(_440_) );
NOR2X1 NOR2X1_41 ( .A(_440_), .B(_439_), .Y(_441_) );
NOR2X1 NOR2X1_42 ( .A(_438_), .B(_441_), .Y(_443_) );
NAND3X1 NAND3X1_57 ( .A(_435_), .B(_437_), .C(_443_), .Y(_444_) );
NOR2X1 NOR2X1_43 ( .A(_433_), .B(_444_), .Y(_445_) );
AOI21X1 AOI21X1_38 ( .A(_386_), .B(_445_), .C(_422_), .Y(_446_) );
INVX1 INVX1_41 ( .A(_338_), .Y(_447_) );
NOR2X1 NOR2X1_44 ( .A(B[7]), .B(A[7]), .Y(_448_) );
OAI21X1 OAI21X1_77 ( .A(_448_), .B(_447_), .C(_445_), .Y(_449_) );
NAND2X1 NAND2X1_45 ( .A(_255_), .B(_421_), .Y(_450_) );
INVX1 INVX1_42 ( .A(_428_), .Y(_451_) );
NOR2X1 NOR2X1_45 ( .A(select[2]), .B(_418_), .Y(_452_) );
INVX1 INVX1_43 ( .A(_452_), .Y(_454_) );
NOR2X1 NOR2X1_46 ( .A(_454_), .B(_266_), .Y(_455_) );
INVX1 INVX1_44 ( .A(_455_), .Y(_456_) );
INVX1 INVX1_45 ( .A(_417_), .Y(_457_) );
NOR2X1 NOR2X1_47 ( .A(_457_), .B(_454_), .Y(_458_) );
NOR2X1 NOR2X1_48 ( .A(select[1]), .B(_244_), .Y(_459_) );
INVX2 INVX2_6 ( .A(_459_), .Y(_460_) );
NOR2X1 NOR2X1_49 ( .A(select[1]), .B(select[0]), .Y(_461_) );
INVX1 INVX1_46 ( .A(_461_), .Y(_462_) );
NOR2X1 NOR2X1_50 ( .A(_222_), .B(_462_), .Y(_463_) );
INVX1 INVX1_47 ( .A(_463_), .Y(_465_) );
OAI21X1 OAI21X1_78 ( .A(_222_), .B(_460_), .C(_465_), .Y(_466_) );
NOR2X1 NOR2X1_51 ( .A(_458_), .B(_466_), .Y(_467_) );
OAI21X1 OAI21X1_79 ( .A(_429_), .B(_467_), .C(_456_), .Y(_468_) );
NOR2X1 NOR2X1_52 ( .A(_222_), .B(_457_), .Y(_469_) );
NOR2X1 NOR2X1_53 ( .A(_462_), .B(_454_), .Y(_470_) );
OAI21X1 OAI21X1_80 ( .A(_469_), .B(_470_), .C(_428_), .Y(_471_) );
INVX1 INVX1_48 ( .A(_421_), .Y(_472_) );
NOR2X1 NOR2X1_54 ( .A(_462_), .B(_472_), .Y(_473_) );
INVX1 INVX1_49 ( .A(_473_), .Y(_474_) );
OAI21X1 OAI21X1_81 ( .A(_472_), .B(_460_), .C(_474_), .Y(_476_) );
NOR2X1 NOR2X1_55 ( .A(select[3]), .B(_419_), .Y(_477_) );
NAND2X1 NAND2X1_46 ( .A(select[0]), .B(_477_), .Y(_478_) );
INVX1 INVX1_50 ( .A(_478_), .Y(_479_) );
AOI22X1 AOI22X1_3 ( .A(A[1]), .B(_479_), .C(_476_), .D(_432_), .Y(_480_) );
INVX1 INVX1_51 ( .A(_429_), .Y(_481_) );
INVX1 INVX1_52 ( .A(_477_), .Y(_482_) );
NOR2X1 NOR2X1_56 ( .A(_457_), .B(_482_), .Y(_483_) );
NOR2X1 NOR2X1_57 ( .A(_454_), .B(_460_), .Y(_484_) );
AOI22X1 AOI22X1_4 ( .A(_483_), .B(A[7]), .C(_481_), .D(_484_), .Y(_485_) );
NAND3X1 NAND3X1_58 ( .A(_471_), .B(_485_), .C(_480_), .Y(_487_) );
AOI21X1 AOI21X1_39 ( .A(_451_), .B(_468_), .C(_487_), .Y(_488_) );
OAI21X1 OAI21X1_82 ( .A(_450_), .B(_449_), .C(_488_), .Y(_489_) );
AOI21X1 AOI21X1_40 ( .A(_416_), .B(_446_), .C(_489_), .Y(_490_) );
OAI21X1 OAI21X1_83 ( .A(_288_), .B(_385_), .C(_490_), .Y(_0__0_) );
XOR2X1 XOR2X1_7 ( .A(_397_), .B(_428_), .Y(_491_) );
NAND2X1 NAND2X1_47 ( .A(_463_), .B(_491_), .Y(_492_) );
OAI21X1 OAI21X1_84 ( .A(_474_), .B(_491_), .C(_492_), .Y(_493_) );
INVX1 INVX1_53 ( .A(_395_), .Y(_494_) );
NOR2X1 NOR2X1_58 ( .A(_494_), .B(_451_), .Y(_495_) );
NAND2X1 NAND2X1_48 ( .A(B[0]), .B(A[1]), .Y(_497_) );
OAI21X1 OAI21X1_85 ( .A(_427_), .B(_387__bF_buf2), .C(_497_), .Y(_498_) );
NAND2X1 NAND2X1_49 ( .A(_498_), .B(_469_), .Y(_499_) );
NOR2X1 NOR2X1_59 ( .A(select[0]), .B(_482_), .Y(_500_) );
NAND2X1 NAND2X1_50 ( .A(A[0]), .B(_500_), .Y(_501_) );
OAI21X1 OAI21X1_86 ( .A(_247_), .B(_478_), .C(_501_), .Y(_502_) );
INVX1 INVX1_54 ( .A(_470_), .Y(_503_) );
OAI21X1 OAI21X1_87 ( .A(B_1_bF_buf0_), .B(A[1]), .C(_484_), .Y(_504_) );
OAI21X1 OAI21X1_88 ( .A(_494_), .B(_503_), .C(_504_), .Y(_505_) );
NOR2X1 NOR2X1_60 ( .A(_502_), .B(_505_), .Y(_506_) );
OAI21X1 OAI21X1_89 ( .A(_495_), .B(_499_), .C(_506_), .Y(_508_) );
NOR2X1 NOR2X1_61 ( .A(_460_), .B(_472_), .Y(_509_) );
INVX1 INVX1_55 ( .A(_509_), .Y(_510_) );
NOR2X1 NOR2X1_62 ( .A(_222_), .B(_460_), .Y(_511_) );
NAND2X1 NAND2X1_51 ( .A(_310_), .B(_397_), .Y(_512_) );
AND2X2 AND2X2_6 ( .A(_400_), .B(_512_), .Y(_513_) );
INVX2 INVX2_7 ( .A(_458_), .Y(_514_) );
OAI21X1 OAI21X1_90 ( .A(_396_), .B(_514_), .C(_456_), .Y(_515_) );
AOI22X1 AOI22X1_5 ( .A(_494_), .B(_515_), .C(_513_), .D(_511_), .Y(_516_) );
OAI21X1 OAI21X1_91 ( .A(_397_), .B(_510_), .C(_516_), .Y(_517_) );
OR2X2 OR2X2_1 ( .A(_517_), .B(_508_), .Y(_519_) );
NOR2X1 NOR2X1_63 ( .A(_493_), .B(_519_), .Y(_520_) );
OAI21X1 OAI21X1_92 ( .A(_288_), .B(_300_), .C(_520_), .Y(_0__1_) );
INVX1 INVX1_56 ( .A(_174_), .Y(_521_) );
OAI21X1 OAI21X1_93 ( .A(_396_), .B(_451_), .C(_494_), .Y(_522_) );
XOR2X1 XOR2X1_8 ( .A(_522_), .B(_438_), .Y(_523_) );
INVX1 INVX1_57 ( .A(_438_), .Y(_524_) );
NAND2X1 NAND2X1_52 ( .A(_211_), .B(_459_), .Y(_525_) );
OAI21X1 OAI21X1_94 ( .A(_525_), .B(_401_), .C(_510_), .Y(_526_) );
AOI22X1 AOI22X1_6 ( .A(_463_), .B(_523_), .C(_526_), .D(_524_), .Y(_527_) );
OAI21X1 OAI21X1_95 ( .A(_474_), .B(_523_), .C(_527_), .Y(_529_) );
NAND2X1 NAND2X1_53 ( .A(A[0]), .B(B_2_bF_buf3_), .Y(_530_) );
NAND2X1 NAND2X1_54 ( .A(B[0]), .B(A[2]), .Y(_531_) );
OAI21X1 OAI21X1_96 ( .A(_387__bF_buf1), .B(_394_), .C(_531_), .Y(_532_) );
NAND2X1 NAND2X1_55 ( .A(A[2]), .B(B_1_bF_buf3_), .Y(_533_) );
OAI21X1 OAI21X1_97 ( .A(_497_), .B(_533_), .C(_532_), .Y(_534_) );
OR2X2 OR2X2_2 ( .A(_534_), .B(_530_), .Y(_535_) );
OAI21X1 OAI21X1_98 ( .A(_427_), .B(_486__bF_buf3), .C(_534_), .Y(_536_) );
AND2X2 AND2X2_7 ( .A(_535_), .B(_536_), .Y(_537_) );
NAND2X1 NAND2X1_56 ( .A(_495_), .B(_537_), .Y(_538_) );
INVX1 INVX1_58 ( .A(_538_), .Y(_540_) );
OAI21X1 OAI21X1_99 ( .A(_495_), .B(_537_), .C(_469_), .Y(_541_) );
NAND2X1 NAND2X1_57 ( .A(_511_), .B(_401_), .Y(_542_) );
OAI21X1 OAI21X1_100 ( .A(_457_), .B(_454_), .C(_542_), .Y(_543_) );
NOR2X1 NOR2X1_64 ( .A(_104_), .B(_478_), .Y(_544_) );
AOI21X1 AOI21X1_41 ( .A(_402_), .B(_470_), .C(_544_), .Y(_545_) );
OAI21X1 OAI21X1_101 ( .A(B_2_bF_buf2_), .B(A[2]), .C(_484_), .Y(_546_) );
INVX1 INVX1_59 ( .A(_402_), .Y(_547_) );
AOI22X1 AOI22X1_7 ( .A(_500_), .B(A[1]), .C(_547_), .D(_455_), .Y(_548_) );
NAND3X1 NAND3X1_59 ( .A(_546_), .B(_545_), .C(_548_), .Y(_549_) );
AOI21X1 AOI21X1_42 ( .A(_543_), .B(_438_), .C(_549_), .Y(_551_) );
OAI21X1 OAI21X1_102 ( .A(_540_), .B(_541_), .C(_551_), .Y(_552_) );
NOR2X1 NOR2X1_65 ( .A(_529_), .B(_552_), .Y(_553_) );
OAI21X1 OAI21X1_103 ( .A(_288_), .B(_521_), .C(_553_), .Y(_0__2_) );
AOI21X1 AOI21X1_43 ( .A(_522_), .B(_438_), .C(_402_), .Y(_554_) );
XOR2X1 XOR2X1_9 ( .A(_554_), .B(_425_), .Y(_555_) );
NAND2X1 NAND2X1_58 ( .A(A[2]), .B(_500_), .Y(_556_) );
OAI21X1 OAI21X1_104 ( .A(_79_), .B(_478_), .C(_556_), .Y(_557_) );
XOR2X1 XOR2X1_10 ( .A(_405_), .B(_426_), .Y(_558_) );
NAND2X1 NAND2X1_59 ( .A(_511_), .B(_558_), .Y(_559_) );
NOR2X1 NOR2X1_66 ( .A(_427_), .B(_431_), .Y(_561_) );
OAI21X1 OAI21X1_105 ( .A(_494_), .B(_531_), .C(_535_), .Y(_562_) );
OAI21X1 OAI21X1_106 ( .A(_299__bF_buf2), .B(_104_), .C(_533_), .Y(_563_) );
NAND2X1 NAND2X1_60 ( .A(A[3]), .B(B_1_bF_buf2_), .Y(_564_) );
OAI21X1 OAI21X1_107 ( .A(_531_), .B(_564_), .C(_563_), .Y(_565_) );
INVX1 INVX1_60 ( .A(_565_), .Y(_566_) );
NAND3X1 NAND3X1_60 ( .A(B_2_bF_buf1_), .B(A[1]), .C(_566_), .Y(_567_) );
OAI21X1 OAI21X1_108 ( .A(_486__bF_buf2), .B(_394_), .C(_565_), .Y(_568_) );
AND2X2 AND2X2_8 ( .A(_567_), .B(_568_), .Y(_569_) );
NAND2X1 NAND2X1_61 ( .A(_562_), .B(_569_), .Y(_570_) );
INVX1 INVX1_61 ( .A(_570_), .Y(_572_) );
NOR2X1 NOR2X1_67 ( .A(_562_), .B(_569_), .Y(_573_) );
NOR2X1 NOR2X1_68 ( .A(_573_), .B(_572_), .Y(_574_) );
XOR2X1 XOR2X1_11 ( .A(_574_), .B(_561_), .Y(_575_) );
OAI21X1 OAI21X1_109 ( .A(_540_), .B(_575_), .C(_469_), .Y(_576_) );
AOI21X1 AOI21X1_44 ( .A(_540_), .B(_575_), .C(_576_), .Y(_577_) );
AOI21X1 AOI21X1_45 ( .A(_92_), .B(_277_), .C(_577_), .Y(_578_) );
NAND2X1 NAND2X1_62 ( .A(_559_), .B(_578_), .Y(_579_) );
OR2X2 OR2X2_3 ( .A(_579_), .B(_557_), .Y(_580_) );
INVX1 INVX1_62 ( .A(_423_), .Y(_581_) );
AOI22X1 AOI22X1_8 ( .A(_455_), .B(_581_), .C(_425_), .D(_458_), .Y(_583_) );
INVX1 INVX1_63 ( .A(_424_), .Y(_584_) );
AOI22X1 AOI22X1_9 ( .A(_470_), .B(_423_), .C(_584_), .D(_484_), .Y(_585_) );
AOI22X1 AOI22X1_10 ( .A(_426_), .B(_509_), .C(_555_), .D(_473_), .Y(_586_) );
NAND3X1 NAND3X1_61 ( .A(_583_), .B(_585_), .C(_586_), .Y(_587_) );
NOR2X1 NOR2X1_69 ( .A(_587_), .B(_580_), .Y(_588_) );
OAI21X1 OAI21X1_110 ( .A(_465_), .B(_555_), .C(_588_), .Y(_0__3_) );
OAI21X1 OAI21X1_111 ( .A(_424_), .B(_554_), .C(_581_), .Y(_589_) );
XOR2X1 XOR2X1_12 ( .A(_589_), .B(_437_), .Y(_590_) );
AOI21X1 AOI21X1_46 ( .A(_407_), .B(_437_), .C(_525_), .Y(_591_) );
OAI21X1 OAI21X1_112 ( .A(_407_), .B(_437_), .C(_591_), .Y(_593_) );
AOI22X1 AOI22X1_11 ( .A(A[5]), .B(_479_), .C(_500_), .D(A[3]), .Y(_594_) );
NAND2X1 NAND2X1_63 ( .A(_540_), .B(_575_), .Y(_595_) );
INVX1 INVX1_64 ( .A(_561_), .Y(_596_) );
OAI21X1 OAI21X1_113 ( .A(_596_), .B(_573_), .C(_570_), .Y(_597_) );
OAI22X1 OAI22X1_2 ( .A(_427_), .B(_376_), .C(_431_), .D(_394_), .Y(_598_) );
NOR2X1 NOR2X1_70 ( .A(_376_), .B(_394_), .Y(_599_) );
INVX1 INVX1_65 ( .A(_599_), .Y(_600_) );
OAI21X1 OAI21X1_114 ( .A(_596_), .B(_600_), .C(_598_), .Y(_601_) );
OAI21X1 OAI21X1_115 ( .A(_107_), .B(_533_), .C(_567_), .Y(_602_) );
OAI21X1 OAI21X1_116 ( .A(_299__bF_buf1), .B(_79_), .C(_564_), .Y(_604_) );
NAND2X1 NAND2X1_64 ( .A(A[4]), .B(B_1_bF_buf1_), .Y(_605_) );
OAI21X1 OAI21X1_117 ( .A(_605_), .B(_107_), .C(_604_), .Y(_606_) );
OAI21X1 OAI21X1_118 ( .A(_486__bF_buf1), .B(_247_), .C(_606_), .Y(_607_) );
OR2X2 OR2X2_4 ( .A(_606_), .B(_547_), .Y(_608_) );
AND2X2 AND2X2_9 ( .A(_608_), .B(_607_), .Y(_609_) );
NAND2X1 NAND2X1_65 ( .A(_602_), .B(_609_), .Y(_610_) );
INVX1 INVX1_66 ( .A(_610_), .Y(_611_) );
NOR2X1 NOR2X1_71 ( .A(_602_), .B(_609_), .Y(_612_) );
NOR2X1 NOR2X1_72 ( .A(_612_), .B(_611_), .Y(_613_) );
XNOR2X1 XNOR2X1_1 ( .A(_613_), .B(_601_), .Y(_615_) );
XNOR2X1 XNOR2X1_2 ( .A(_615_), .B(_597_), .Y(_616_) );
NOR2X1 NOR2X1_73 ( .A(_595_), .B(_616_), .Y(_617_) );
INVX1 INVX1_67 ( .A(_617_), .Y(_618_) );
INVX1 INVX1_68 ( .A(_469_), .Y(_619_) );
AOI21X1 AOI21X1_47 ( .A(_616_), .B(_595_), .C(_619_), .Y(_620_) );
AOI22X1 AOI22X1_12 ( .A(_618_), .B(_620_), .C(_45_), .D(_277_), .Y(_621_) );
NAND3X1 NAND3X1_62 ( .A(_593_), .B(_594_), .C(_621_), .Y(_622_) );
INVX1 INVX1_69 ( .A(_410_), .Y(_623_) );
AOI22X1 AOI22X1_13 ( .A(_470_), .B(_408_), .C(_623_), .D(_484_), .Y(_624_) );
OAI21X1 OAI21X1_119 ( .A(_410_), .B(_514_), .C(_456_), .Y(_626_) );
OAI21X1 OAI21X1_120 ( .A(_376_), .B(_79_), .C(_626_), .Y(_627_) );
AOI22X1 AOI22X1_14 ( .A(_437_), .B(_509_), .C(_590_), .D(_473_), .Y(_628_) );
NAND3X1 NAND3X1_63 ( .A(_624_), .B(_627_), .C(_628_), .Y(_629_) );
NOR2X1 NOR2X1_74 ( .A(_629_), .B(_622_), .Y(_630_) );
OAI21X1 OAI21X1_121 ( .A(_465_), .B(_590_), .C(_630_), .Y(_0__4_) );
NAND2X1 NAND2X1_66 ( .A(_597_), .B(_615_), .Y(_631_) );
INVX1 INVX1_70 ( .A(_631_), .Y(_632_) );
NOR2X1 NOR2X1_75 ( .A(_596_), .B(_600_), .Y(_633_) );
OAI21X1 OAI21X1_122 ( .A(_601_), .B(_612_), .C(_610_), .Y(_634_) );
NOR2X1 NOR2X1_76 ( .A(_427_), .B(_409_), .Y(_636_) );
NAND2X1 NAND2X1_67 ( .A(B[3]), .B(A[2]), .Y(_637_) );
XNOR2X1 XNOR2X1_3 ( .A(_599_), .B(_637_), .Y(_638_) );
XOR2X1 XOR2X1_13 ( .A(_638_), .B(_636_), .Y(_639_) );
OAI21X1 OAI21X1_123 ( .A(_107_), .B(_605_), .C(_608_), .Y(_640_) );
XOR2X1 XOR2X1_14 ( .A(_35_), .B(_605_), .Y(_641_) );
INVX1 INVX1_71 ( .A(_641_), .Y(_642_) );
NAND3X1 NAND3X1_64 ( .A(A[3]), .B(B_2_bF_buf0_), .C(_642_), .Y(_643_) );
OAI21X1 OAI21X1_124 ( .A(_104_), .B(_486__bF_buf0), .C(_641_), .Y(_644_) );
AND2X2 AND2X2_10 ( .A(_643_), .B(_644_), .Y(_645_) );
XOR2X1 XOR2X1_15 ( .A(_645_), .B(_640_), .Y(_647_) );
XOR2X1 XOR2X1_16 ( .A(_647_), .B(_639_), .Y(_648_) );
NAND2X1 NAND2X1_68 ( .A(_634_), .B(_648_), .Y(_649_) );
INVX1 INVX1_72 ( .A(_649_), .Y(_650_) );
NOR2X1 NOR2X1_77 ( .A(_634_), .B(_648_), .Y(_651_) );
NOR2X1 NOR2X1_78 ( .A(_651_), .B(_650_), .Y(_652_) );
XOR2X1 XOR2X1_17 ( .A(_652_), .B(_633_), .Y(_653_) );
NAND2X1 NAND2X1_69 ( .A(_632_), .B(_653_), .Y(_654_) );
INVX1 INVX1_73 ( .A(_654_), .Y(_655_) );
NOR2X1 NOR2X1_79 ( .A(_632_), .B(_653_), .Y(_656_) );
OAI21X1 OAI21X1_125 ( .A(_656_), .B(_655_), .C(_618_), .Y(_658_) );
NAND2X1 NAND2X1_70 ( .A(_617_), .B(_653_), .Y(_659_) );
INVX1 INVX1_74 ( .A(_659_), .Y(_660_) );
NOR2X1 NOR2X1_80 ( .A(_619_), .B(_660_), .Y(_661_) );
AND2X2 AND2X2_11 ( .A(_412_), .B(_441_), .Y(_662_) );
NOR2X1 NOR2X1_81 ( .A(_441_), .B(_412_), .Y(_663_) );
OAI21X1 OAI21X1_126 ( .A(_663_), .B(_662_), .C(_511_), .Y(_664_) );
NAND2X1 NAND2X1_71 ( .A(_436_), .B(_589_), .Y(_665_) );
OAI21X1 OAI21X1_127 ( .A(_376_), .B(_79_), .C(_665_), .Y(_666_) );
XOR2X1 XOR2X1_18 ( .A(_666_), .B(_441_), .Y(_667_) );
NAND2X1 NAND2X1_72 ( .A(_463_), .B(_667_), .Y(_669_) );
NOR2X1 NOR2X1_82 ( .A(_474_), .B(_667_), .Y(_670_) );
INVX1 INVX1_75 ( .A(_439_), .Y(_671_) );
OAI21X1 OAI21X1_128 ( .A(_440_), .B(_514_), .C(_456_), .Y(_672_) );
INVX1 INVX1_76 ( .A(_440_), .Y(_673_) );
AOI22X1 AOI22X1_15 ( .A(_500_), .B(A[4]), .C(_673_), .D(_484_), .Y(_674_) );
OAI21X1 OAI21X1_129 ( .A(_389_), .B(_478_), .C(_674_), .Y(_675_) );
INVX1 INVX1_77 ( .A(_675_), .Y(_676_) );
OAI21X1 OAI21X1_130 ( .A(_671_), .B(_503_), .C(_676_), .Y(_677_) );
AOI21X1 AOI21X1_48 ( .A(_671_), .B(_672_), .C(_677_), .Y(_678_) );
OAI21X1 OAI21X1_131 ( .A(_441_), .B(_510_), .C(_678_), .Y(_680_) );
NOR2X1 NOR2X1_83 ( .A(_680_), .B(_670_), .Y(_681_) );
NAND3X1 NAND3X1_65 ( .A(_669_), .B(_681_), .C(_664_), .Y(_682_) );
AOI21X1 AOI21X1_49 ( .A(_661_), .B(_658_), .C(_682_), .Y(_683_) );
OAI21X1 OAI21X1_132 ( .A(_288_), .B(_50_), .C(_683_), .Y(_0__5_) );
INVX1 INVX1_78 ( .A(_633_), .Y(_684_) );
OAI21X1 OAI21X1_133 ( .A(_684_), .B(_651_), .C(_649_), .Y(_685_) );
NOR2X1 NOR2X1_84 ( .A(_427_), .B(_398_), .Y(_686_) );
NAND2X1 NAND2X1_73 ( .A(_636_), .B(_638_), .Y(_687_) );
OAI21X1 OAI21X1_134 ( .A(_600_), .B(_637_), .C(_687_), .Y(_688_) );
XOR2X1 XOR2X1_19 ( .A(_688_), .B(_686_), .Y(_690_) );
NAND2X1 NAND2X1_74 ( .A(_640_), .B(_645_), .Y(_691_) );
NAND2X1 NAND2X1_75 ( .A(_639_), .B(_647_), .Y(_692_) );
NAND2X1 NAND2X1_76 ( .A(_691_), .B(_692_), .Y(_693_) );
NAND2X1 NAND2X1_77 ( .A(B[4]), .B(A[2]), .Y(_694_) );
OAI21X1 OAI21X1_135 ( .A(_431_), .B(_104_), .C(_694_), .Y(_695_) );
NAND2X1 NAND2X1_78 ( .A(B[4]), .B(A[3]), .Y(_696_) );
OAI21X1 OAI21X1_136 ( .A(_637_), .B(_696_), .C(_695_), .Y(_697_) );
INVX1 INVX1_79 ( .A(_697_), .Y(_698_) );
NAND3X1 NAND3X1_66 ( .A(B[5]), .B(A[1]), .C(_698_), .Y(_699_) );
OAI21X1 OAI21X1_137 ( .A(_409_), .B(_394_), .C(_697_), .Y(_701_) );
NAND2X1 NAND2X1_79 ( .A(_701_), .B(_699_), .Y(_702_) );
OAI21X1 OAI21X1_138 ( .A(_36_), .B(_605_), .C(_643_), .Y(_703_) );
NAND2X1 NAND2X1_80 ( .A(A[4]), .B(B_2_bF_buf3_), .Y(_704_) );
OAI22X1 OAI22X1_3 ( .A(_299__bF_buf0), .B(_389_), .C(_21_), .D(_387__bF_buf0), .Y(_705_) );
NOR2X1 NOR2X1_85 ( .A(_389_), .B(_387__bF_buf3), .Y(_706_) );
INVX1 INVX1_80 ( .A(_706_), .Y(_707_) );
OAI21X1 OAI21X1_139 ( .A(_36_), .B(_707_), .C(_705_), .Y(_708_) );
OR2X2 OR2X2_5 ( .A(_708_), .B(_704_), .Y(_709_) );
OAI21X1 OAI21X1_140 ( .A(_79_), .B(_486__bF_buf3), .C(_708_), .Y(_710_) );
AND2X2 AND2X2_12 ( .A(_709_), .B(_710_), .Y(_712_) );
NAND2X1 NAND2X1_81 ( .A(_703_), .B(_712_), .Y(_713_) );
INVX1 INVX1_81 ( .A(_713_), .Y(_714_) );
NOR2X1 NOR2X1_86 ( .A(_703_), .B(_712_), .Y(_715_) );
NOR2X1 NOR2X1_87 ( .A(_715_), .B(_714_), .Y(_716_) );
XNOR2X1 XNOR2X1_4 ( .A(_716_), .B(_702_), .Y(_717_) );
NAND2X1 NAND2X1_82 ( .A(_693_), .B(_717_), .Y(_718_) );
INVX1 INVX1_82 ( .A(_718_), .Y(_719_) );
NOR2X1 NOR2X1_88 ( .A(_693_), .B(_717_), .Y(_720_) );
NOR2X1 NOR2X1_89 ( .A(_720_), .B(_719_), .Y(_721_) );
XOR2X1 XOR2X1_20 ( .A(_721_), .B(_690_), .Y(_723_) );
XNOR2X1 XNOR2X1_5 ( .A(_723_), .B(_685_), .Y(_724_) );
OR2X2 OR2X2_6 ( .A(_724_), .B(_654_), .Y(_725_) );
NAND2X1 NAND2X1_83 ( .A(_654_), .B(_724_), .Y(_726_) );
AND2X2 AND2X2_13 ( .A(_725_), .B(_726_), .Y(_727_) );
OAI21X1 OAI21X1_141 ( .A(_660_), .B(_727_), .C(_469_), .Y(_728_) );
AOI21X1 AOI21X1_50 ( .A(_660_), .B(_727_), .C(_728_), .Y(_729_) );
INVX1 INVX1_83 ( .A(_666_), .Y(_730_) );
OAI21X1 OAI21X1_142 ( .A(_440_), .B(_730_), .C(_671_), .Y(_731_) );
XOR2X1 XOR2X1_21 ( .A(_731_), .B(_434_), .Y(_732_) );
OAI21X1 OAI21X1_143 ( .A(B[6]), .B(A[6]), .C(_484_), .Y(_734_) );
OAI21X1 OAI21X1_144 ( .A(_392_), .B(_456_), .C(_734_), .Y(_735_) );
INVX1 INVX1_84 ( .A(A[7]), .Y(_736_) );
OAI22X1 OAI22X1_4 ( .A(_736_), .B(_478_), .C(_435_), .D(_514_), .Y(_737_) );
OR2X2 OR2X2_7 ( .A(_737_), .B(_735_), .Y(_738_) );
AOI22X1 AOI22X1_16 ( .A(_500_), .B(A[5]), .C(_392_), .D(_470_), .Y(_739_) );
OAI21X1 OAI21X1_145 ( .A(_434_), .B(_510_), .C(_739_), .Y(_740_) );
NOR2X1 NOR2X1_90 ( .A(_740_), .B(_738_), .Y(_741_) );
OAI21X1 OAI21X1_146 ( .A(_288_), .B(_711_), .C(_741_), .Y(_742_) );
NOR2X1 NOR2X1_91 ( .A(_435_), .B(_414_), .Y(_743_) );
NAND2X1 NAND2X1_84 ( .A(_511_), .B(_415_), .Y(_745_) );
NAND2X1 NAND2X1_85 ( .A(_463_), .B(_732_), .Y(_746_) );
OAI21X1 OAI21X1_147 ( .A(_743_), .B(_745_), .C(_746_), .Y(_747_) );
NOR2X1 NOR2X1_92 ( .A(_742_), .B(_747_), .Y(_748_) );
OAI21X1 OAI21X1_148 ( .A(_474_), .B(_732_), .C(_748_), .Y(_749_) );
OR2X2 OR2X2_8 ( .A(_729_), .B(_749_), .Y(_0__6_) );
AND2X2 AND2X2_14 ( .A(_507_), .B(_453_), .Y(_750_) );
NAND3X1 NAND3X1_67 ( .A(A[0]), .B(_477_), .C(_255_), .Y(_751_) );
NAND2X1 NAND2X1_86 ( .A(A[6]), .B(_500_), .Y(_752_) );
OAI21X1 OAI21X1_149 ( .A(B[7]), .B(A[7]), .C(_484_), .Y(_753_) );
NAND3X1 NAND3X1_68 ( .A(_751_), .B(_752_), .C(_753_), .Y(_755_) );
AOI21X1 AOI21X1_51 ( .A(_277_), .B(_750_), .C(_755_), .Y(_756_) );
NAND2X1 NAND2X1_87 ( .A(_470_), .B(_447_), .Y(_757_) );
AND2X2 AND2X2_15 ( .A(_757_), .B(_756_), .Y(_758_) );
INVX1 INVX1_85 ( .A(_727_), .Y(_759_) );
OAI21X1 OAI21X1_150 ( .A(_659_), .B(_759_), .C(_725_), .Y(_760_) );
AOI21X1 AOI21X1_52 ( .A(_721_), .B(_690_), .C(_719_), .Y(_761_) );
OAI21X1 OAI21X1_151 ( .A(_36_), .B(_707_), .C(_709_), .Y(_762_) );
NOR2X1 NOR2X1_93 ( .A(_21_), .B(_486__bF_buf2), .Y(_763_) );
NOR2X1 NOR2X1_94 ( .A(_299__bF_buf3), .B(_736_), .Y(_764_) );
XNOR2X1 XNOR2X1_6 ( .A(_764_), .B(_706_), .Y(_766_) );
XNOR2X1 XNOR2X1_7 ( .A(_766_), .B(_763_), .Y(_767_) );
XNOR2X1 XNOR2X1_8 ( .A(_762_), .B(_767_), .Y(_768_) );
NOR2X1 NOR2X1_95 ( .A(_409_), .B(_247_), .Y(_769_) );
NAND2X1 NAND2X1_88 ( .A(A[4]), .B(B[3]), .Y(_770_) );
XNOR2X1 XNOR2X1_9 ( .A(_696_), .B(_770_), .Y(_771_) );
XOR2X1 XOR2X1_22 ( .A(_771_), .B(_769_), .Y(_772_) );
NAND2X1 NAND2X1_89 ( .A(A[0]), .B(B[7]), .Y(_773_) );
NAND2X1 NAND2X1_90 ( .A(B[6]), .B(A[1]), .Y(_774_) );
XNOR2X1 XNOR2X1_10 ( .A(_773_), .B(_774_), .Y(_775_) );
XOR2X1 XOR2X1_23 ( .A(_772_), .B(_775_), .Y(_777_) );
XOR2X1 XOR2X1_24 ( .A(_768_), .B(_777_), .Y(_778_) );
OAI21X1 OAI21X1_152 ( .A(_581_), .B(_694_), .C(_699_), .Y(_779_) );
OAI21X1 OAI21X1_153 ( .A(_702_), .B(_715_), .C(_713_), .Y(_780_) );
XOR2X1 XOR2X1_25 ( .A(_780_), .B(_779_), .Y(_781_) );
XOR2X1 XOR2X1_26 ( .A(_781_), .B(_778_), .Y(_782_) );
XOR2X1 XOR2X1_27 ( .A(_761_), .B(_782_), .Y(_783_) );
NAND2X1 NAND2X1_91 ( .A(_686_), .B(_688_), .Y(_784_) );
NAND2X1 NAND2X1_92 ( .A(_685_), .B(_723_), .Y(_785_) );
XOR2X1 XOR2X1_28 ( .A(_785_), .B(_784_), .Y(_786_) );
XOR2X1 XOR2X1_29 ( .A(_786_), .B(_783_), .Y(_788_) );
OAI21X1 OAI21X1_154 ( .A(_788_), .B(_760_), .C(_469_), .Y(_789_) );
AOI21X1 AOI21X1_53 ( .A(_760_), .B(_788_), .C(_789_), .Y(_790_) );
AOI21X1 AOI21X1_54 ( .A(_338_), .B(_455_), .C(_790_), .Y(_791_) );
AND2X2 AND2X2_16 ( .A(_758_), .B(_791_), .Y(_792_) );
OAI21X1 OAI21X1_155 ( .A(B[6]), .B(_389_), .C(_415_), .Y(_793_) );
INVX1 INVX1_86 ( .A(_793_), .Y(_794_) );
OAI21X1 OAI21X1_156 ( .A(_525_), .B(_794_), .C(_514_), .Y(_795_) );
AOI21X1 AOI21X1_55 ( .A(_794_), .B(_511_), .C(_509_), .Y(_796_) );
OAI21X1 OAI21X1_157 ( .A(_448_), .B(_447_), .C(_796_), .Y(_797_) );
OAI21X1 OAI21X1_158 ( .A(_386_), .B(_795_), .C(_797_), .Y(_799_) );
AOI21X1 AOI21X1_56 ( .A(_731_), .B(_434_), .C(_392_), .Y(_800_) );
NOR2X1 NOR2X1_96 ( .A(_800_), .B(_386_), .Y(_801_) );
INVX1 INVX1_87 ( .A(_801_), .Y(_802_) );
OAI21X1 OAI21X1_159 ( .A(_448_), .B(_447_), .C(_800_), .Y(_803_) );
NAND2X1 NAND2X1_93 ( .A(_803_), .B(_802_), .Y(_804_) );
MUX2X1 MUX2X1_1 ( .A(_473_), .B(_463_), .S(_804_), .Y(_805_) );
NAND3X1 NAND3X1_69 ( .A(_792_), .B(_799_), .C(_805_), .Y(_0__7_) );
OAI21X1 OAI21X1_160 ( .A(_448_), .B(_800_), .C(_338_), .Y(_822_) );
BUFX2 BUFX2_20 ( .A(_821__0_), .Y(ALU_out[0]) );
BUFX2 BUFX2_21 ( .A(_821__1_), .Y(ALU_out[1]) );
BUFX2 BUFX2_22 ( .A(_821__2_), .Y(ALU_out[2]) );
BUFX2 BUFX2_23 ( .A(_821__3_), .Y(ALU_out[3]) );
BUFX2 BUFX2_24 ( .A(_821__4_), .Y(ALU_out[4]) );
BUFX2 BUFX2_25 ( .A(_821__5_), .Y(ALU_out[5]) );
BUFX2 BUFX2_26 ( .A(_821__6_), .Y(ALU_out[6]) );
BUFX2 BUFX2_27 ( .A(_821__7_), .Y(ALU_out[7]) );
BUFX2 BUFX2_28 ( .A(_822_), .Y(Carry_out) );
DFFPOSX1 DFFPOSX1_1 ( .CLK(clk), .D(_0__0_), .Q(_821__0_) );
DFFPOSX1 DFFPOSX1_2 ( .CLK(clk), .D(_0__1_), .Q(_821__1_) );
DFFPOSX1 DFFPOSX1_3 ( .CLK(clk), .D(_0__2_), .Q(_821__2_) );
DFFPOSX1 DFFPOSX1_4 ( .CLK(clk), .D(_0__3_), .Q(_821__3_) );
DFFPOSX1 DFFPOSX1_5 ( .CLK(clk), .D(_0__4_), .Q(_821__4_) );
DFFPOSX1 DFFPOSX1_6 ( .CLK(clk), .D(_0__5_), .Q(_821__5_) );
DFFPOSX1 DFFPOSX1_7 ( .CLK(clk), .D(_0__6_), .Q(_821__6_) );
DFFPOSX1 DFFPOSX1_8 ( .CLK(clk), .D(_0__7_), .Q(_821__7_) );
NOR2X1 NOR2X1_97 ( .A(select[3]), .B(select[2]), .Y(_211_) );
INVX1 INVX1_88 ( .A(_211_), .Y(_222_) );
INVX1 INVX1_89 ( .A(select[1]), .Y(_233_) );
INVX1 INVX1_90 ( .A(select[0]), .Y(_244_) );
NOR2X1 NOR2X1_98 ( .A(_233_), .B(_244_), .Y(_255_) );
INVX1 INVX1_91 ( .A(_255_), .Y(_266_) );
NOR2X1 NOR2X1_99 ( .A(_222_), .B(_266_), .Y(_277_) );
INVX2 INVX2_8 ( .A(_277_), .Y(_288_) );
INVX4 INVX4_1 ( .A(B[0]), .Y(_299_) );
NOR2X1 NOR2X1_100 ( .A(A[0]), .B(_299__bF_buf2), .Y(_310_) );
NAND2X1 NAND2X1_94 ( .A(B_1_bF_buf0_), .B(_310_), .Y(_321_) );
NOR2X1 NOR2X1_101 ( .A(B[7]), .B(B[6]), .Y(_332_) );
INVX4 INVX4_2 ( .A(_332_), .Y(_343_) );
NOR2X1 NOR2X1_102 ( .A(B[5]), .B(_343_), .Y(_354_) );
INVX4 INVX4_3 ( .A(_354_), .Y(_365_) );
INVX4 INVX4_4 ( .A(B[4]), .Y(_376_) );
INVX4 INVX4_5 ( .A(B_1_bF_buf3_), .Y(_387_) );
INVX1 INVX1_92 ( .A(B[6]), .Y(_398_) );
INVX2 INVX2_9 ( .A(B[5]), .Y(_409_) );
NAND2X1 NAND2X1_95 ( .A(_398_), .B(_409_), .Y(_420_) );
INVX4 INVX4_6 ( .A(B[3]), .Y(_431_) );
NAND2X1 NAND2X1_96 ( .A(_376_), .B(_431_), .Y(_442_) );
NOR2X1 NOR2X1_103 ( .A(_420_), .B(_442_), .Y(_453_) );
INVX2 INVX2_10 ( .A(B[7]), .Y(_464_) );
NAND2X1 NAND2X1_97 ( .A(_464_), .B(_387__bF_buf2), .Y(_475_) );
INVX4 INVX4_7 ( .A(B_2_bF_buf2_), .Y(_486_) );
OAI21X1 OAI21X1_161 ( .A(A[7]), .B(_299__bF_buf1), .C(_486__bF_buf1), .Y(_496_) );
NOR2X1 NOR2X1_104 ( .A(_475_), .B(_496_), .Y(_507_) );
NAND3X1 NAND3X1_70 ( .A(B[0]), .B(_453_), .C(_507_), .Y(_518_) );
NAND3X1 NAND3X1_71 ( .A(A[7]), .B(_387__bF_buf1), .C(_518_), .Y(_528_) );
NOR2X1 NOR2X1_105 ( .A(A[7]), .B(_387__bF_buf0), .Y(_539_) );
INVX1 INVX1_93 ( .A(_539_), .Y(_550_) );
NOR2X1 NOR2X1_106 ( .A(A[6]), .B(_299__bF_buf0), .Y(_560_) );
INVX1 INVX1_94 ( .A(_560_), .Y(_571_) );
NAND3X1 NAND3X1_72 ( .A(_550_), .B(_571_), .C(_528_), .Y(_582_) );
NOR2X1 NOR2X1_107 ( .A(B[5]), .B(B[4]), .Y(_592_) );
NOR2X1 NOR2X1_108 ( .A(B[3]), .B(B_2_bF_buf1_), .Y(_603_) );
NAND3X1 NAND3X1_73 ( .A(_332_), .B(_592_), .C(_603_), .Y(_614_) );
AOI21X1 AOI21X1_57 ( .A(_582_), .B(_528_), .C(_614_), .Y(_625_) );
OAI21X1 OAI21X1_162 ( .A(A[7]), .B(_387__bF_buf3), .C(_528_), .Y(_635_) );
NAND2X1 NAND2X1_98 ( .A(_560_), .B(_635_), .Y(_646_) );
NAND3X1 NAND3X1_74 ( .A(_582_), .B(_646_), .C(_625_), .Y(_657_) );
INVX2 INVX2_11 ( .A(_657_), .Y(_668_) );
NOR2X1 NOR2X1_109 ( .A(B[4]), .B(_365_), .Y(_679_) );
INVX1 INVX1_95 ( .A(_614_), .Y(_689_) );
OAI21X1 OAI21X1_163 ( .A(_539_), .B(_560_), .C(_528_), .Y(_700_) );
NAND2X1 NAND2X1_99 ( .A(_689_), .B(_700_), .Y(_711_) );
NAND3X1 NAND3X1_75 ( .A(A[7]), .B(_518_), .C(_711_), .Y(_722_) );
NAND3X1 NAND3X1_76 ( .A(B[0]), .B(_689_), .C(_700_), .Y(_733_) );
NAND3X1 NAND3X1_77 ( .A(A[6]), .B(_387__bF_buf2), .C(_733_), .Y(_744_) );
NAND2X1 NAND2X1_100 ( .A(A[6]), .B(_733_), .Y(_754_) );
NAND2X1 NAND2X1_101 ( .A(B_1_bF_buf2_), .B(_754_), .Y(_765_) );
NOR2X1 NOR2X1_110 ( .A(A[5]), .B(_299__bF_buf3), .Y(_776_) );
INVX1 INVX1_96 ( .A(_776_), .Y(_787_) );
NAND3X1 NAND3X1_78 ( .A(_744_), .B(_787_), .C(_765_), .Y(_798_) );
NAND3X1 NAND3X1_79 ( .A(B_2_bF_buf0_), .B(_744_), .C(_798_), .Y(_806_) );
AOI21X1 AOI21X1_58 ( .A(_733_), .B(A[6]), .C(_387__bF_buf1), .Y(_807_) );
OAI21X1 OAI21X1_164 ( .A(_776_), .B(_807_), .C(_744_), .Y(_808_) );
NAND2X1 NAND2X1_102 ( .A(_431_), .B(_679_), .Y(_809_) );
AOI21X1 AOI21X1_59 ( .A(_808_), .B(_486__bF_buf0), .C(_809_), .Y(_810_) );
AOI22X1 AOI22X1_17 ( .A(_657_), .B(_722_), .C(_806_), .D(_810_), .Y(_811_) );
INVX1 INVX1_97 ( .A(_811_), .Y(_812_) );
NAND2X1 NAND2X1_103 ( .A(_431_), .B(_811_), .Y(_813_) );
INVX1 INVX1_98 ( .A(_813_), .Y(_814_) );
INVX1 INVX1_99 ( .A(_754_), .Y(_815_) );
AOI21X1 AOI21X1_60 ( .A(_657_), .B(_722_), .C(B_2_bF_buf3_), .Y(_816_) );
NAND3X1 NAND3X1_80 ( .A(B_2_bF_buf2_), .B(_722_), .C(_657_), .Y(_817_) );
AOI21X1 AOI21X1_61 ( .A(_808_), .B(_817_), .C(_816_), .Y(_818_) );
OAI21X1 OAI21X1_165 ( .A(_809_), .B(_818_), .C(_815_), .Y(_819_) );
INVX1 INVX1_100 ( .A(_809_), .Y(_820_) );
NAND2X1 NAND2X1_104 ( .A(_722_), .B(_657_), .Y(_1_) );
NAND2X1 NAND2X1_105 ( .A(_486__bF_buf3), .B(_1_), .Y(_2_) );
NAND2X1 NAND2X1_106 ( .A(_817_), .B(_808_), .Y(_3_) );
NAND2X1 NAND2X1_107 ( .A(_2_), .B(_3_), .Y(_4_) );
INVX1 INVX1_101 ( .A(_744_), .Y(_5_) );
OAI21X1 OAI21X1_166 ( .A(_807_), .B(_5_), .C(_776_), .Y(_6_) );
AND2X2 AND2X2_17 ( .A(_6_), .B(_798_), .Y(_7_) );
NAND3X1 NAND3X1_81 ( .A(_820_), .B(_4_), .C(_7_), .Y(_8_) );
AOI21X1 AOI21X1_62 ( .A(_8_), .B(_819_), .C(B_2_bF_buf1_), .Y(_9_) );
XOR2X1 XOR2X1_30 ( .A(_811_), .B(_431_), .Y(_10_) );
AOI21X1 AOI21X1_63 ( .A(_10_), .B(_9_), .C(_814_), .Y(_11_) );
NAND2X1 NAND2X1_108 ( .A(_798_), .B(_6_), .Y(_12_) );
NAND3X1 NAND3X1_82 ( .A(_820_), .B(_12_), .C(_4_), .Y(_13_) );
OAI21X1 OAI21X1_167 ( .A(_809_), .B(_818_), .C(_754_), .Y(_14_) );
NAND3X1 NAND3X1_83 ( .A(_486__bF_buf2), .B(_14_), .C(_13_), .Y(_15_) );
NAND3X1 NAND3X1_84 ( .A(B_2_bF_buf0_), .B(_819_), .C(_8_), .Y(_16_) );
NAND3X1 NAND3X1_85 ( .A(_15_), .B(_16_), .C(_10_), .Y(_17_) );
NOR2X1 NOR2X1_111 ( .A(_299__bF_buf2), .B(_809_), .Y(_18_) );
INVX1 INVX1_102 ( .A(_18_), .Y(_19_) );
OAI21X1 OAI21X1_168 ( .A(_19_), .B(_818_), .C(A[5]), .Y(_20_) );
INVX2 INVX2_12 ( .A(A[5]), .Y(_21_) );
NAND3X1 NAND3X1_86 ( .A(_21_), .B(_18_), .C(_4_), .Y(_22_) );
AOI21X1 AOI21X1_64 ( .A(_22_), .B(_20_), .C(B_1_bF_buf1_), .Y(_23_) );
NAND3X1 NAND3X1_87 ( .A(B_1_bF_buf0_), .B(_20_), .C(_22_), .Y(_24_) );
NOR2X1 NOR2X1_112 ( .A(A[4]), .B(_299__bF_buf1), .Y(_25_) );
INVX1 INVX1_103 ( .A(_25_), .Y(_26_) );
AOI21X1 AOI21X1_65 ( .A(_24_), .B(_26_), .C(_23_), .Y(_27_) );
OAI21X1 OAI21X1_169 ( .A(_27_), .B(_17_), .C(_11_), .Y(_28_) );
AOI21X1 AOI21X1_66 ( .A(_28_), .B(_679_), .C(_812_), .Y(_29_) );
OAI21X1 OAI21X1_170 ( .A(_668_), .B(_29_), .C(_376_), .Y(_30_) );
NOR3X1 NOR3X1_1 ( .A(_376_), .B(_668_), .C(_29_), .Y(_31_) );
INVX2 INVX2_13 ( .A(_679_), .Y(_32_) );
AND2X2 AND2X2_18 ( .A(_16_), .B(_15_), .Y(_33_) );
NAND2X1 NAND2X1_109 ( .A(_299__bF_buf0), .B(_21_), .Y(_34_) );
NOR2X1 NOR2X1_113 ( .A(_299__bF_buf3), .B(_21_), .Y(_35_) );
INVX1 INVX1_104 ( .A(_35_), .Y(_36_) );
AND2X2 AND2X2_19 ( .A(_36_), .B(_34_), .Y(_37_) );
INVX1 INVX1_105 ( .A(_37_), .Y(_38_) );
NAND3X1 NAND3X1_88 ( .A(_820_), .B(_38_), .C(_4_), .Y(_39_) );
OAI21X1 OAI21X1_171 ( .A(_809_), .B(_818_), .C(_21_), .Y(_40_) );
NAND3X1 NAND3X1_89 ( .A(_387__bF_buf0), .B(_40_), .C(_39_), .Y(_41_) );
AOI21X1 AOI21X1_67 ( .A(_39_), .B(_40_), .C(_387__bF_buf3), .Y(_42_) );
OAI21X1 OAI21X1_172 ( .A(_25_), .B(_42_), .C(_41_), .Y(_43_) );
NAND3X1 NAND3X1_90 ( .A(_10_), .B(_33_), .C(_43_), .Y(_44_) );
AOI21X1 AOI21X1_68 ( .A(_44_), .B(_11_), .C(_32_), .Y(_45_) );
NAND2X1 NAND2X1_110 ( .A(_15_), .B(_16_), .Y(_46_) );
NOR2X1 NOR2X1_114 ( .A(_46_), .B(_27_), .Y(_47_) );
NOR2X1 NOR2X1_115 ( .A(_33_), .B(_43_), .Y(_48_) );
OAI21X1 OAI21X1_173 ( .A(_47_), .B(_48_), .C(_45_), .Y(_49_) );
NAND2X1 NAND2X1_111 ( .A(_820_), .B(_4_), .Y(_50_) );
OAI21X1 OAI21X1_174 ( .A(_12_), .B(_50_), .C(_819_), .Y(_51_) );
INVX1 INVX1_106 ( .A(_51_), .Y(_52_) );
XOR2X1 XOR2X1_31 ( .A(_811_), .B(B[3]), .Y(_53_) );
OAI21X1 OAI21X1_175 ( .A(_15_), .B(_53_), .C(_813_), .Y(_54_) );
NOR2X1 NOR2X1_116 ( .A(_53_), .B(_46_), .Y(_55_) );
AOI21X1 AOI21X1_69 ( .A(_55_), .B(_43_), .C(_54_), .Y(_56_) );
OAI21X1 OAI21X1_176 ( .A(_32_), .B(_56_), .C(_52_), .Y(_57_) );
NAND3X1 NAND3X1_91 ( .A(_431_), .B(_57_), .C(_49_), .Y(_58_) );
OAI21X1 OAI21X1_177 ( .A(_58_), .B(_31_), .C(_30_), .Y(_59_) );
INVX1 INVX1_107 ( .A(_59_), .Y(_60_) );
OAI21X1 OAI21X1_178 ( .A(_32_), .B(_56_), .C(_811_), .Y(_61_) );
NAND3X1 NAND3X1_92 ( .A(_376_), .B(_657_), .C(_61_), .Y(_62_) );
OAI21X1 OAI21X1_179 ( .A(_668_), .B(_29_), .C(B[4]), .Y(_63_) );
XNOR2X1 XNOR2X1_11 ( .A(_43_), .B(_46_), .Y(_64_) );
NAND2X1 NAND2X1_112 ( .A(_64_), .B(_45_), .Y(_65_) );
OAI21X1 OAI21X1_180 ( .A(_32_), .B(_56_), .C(_51_), .Y(_66_) );
NAND3X1 NAND3X1_93 ( .A(_431_), .B(_65_), .C(_66_), .Y(_67_) );
NAND3X1 NAND3X1_94 ( .A(B[3]), .B(_57_), .C(_49_), .Y(_68_) );
AOI22X1 AOI22X1_18 ( .A(_62_), .B(_63_), .C(_67_), .D(_68_), .Y(_69_) );
NAND3X1 NAND3X1_95 ( .A(_26_), .B(_41_), .C(_24_), .Y(_70_) );
OAI21X1 OAI21X1_181 ( .A(_23_), .B(_42_), .C(_25_), .Y(_71_) );
NAND2X1 NAND2X1_113 ( .A(_70_), .B(_71_), .Y(_72_) );
NAND2X1 NAND2X1_114 ( .A(_72_), .B(_45_), .Y(_73_) );
OAI21X1 OAI21X1_182 ( .A(_37_), .B(_50_), .C(_40_), .Y(_74_) );
OAI21X1 OAI21X1_183 ( .A(_32_), .B(_56_), .C(_74_), .Y(_75_) );
AOI21X1 AOI21X1_70 ( .A(_75_), .B(_73_), .C(_486__bF_buf1), .Y(_76_) );
INVX1 INVX1_108 ( .A(_76_), .Y(_77_) );
NAND3X1 NAND3X1_96 ( .A(_486__bF_buf0), .B(_73_), .C(_75_), .Y(_78_) );
INVX2 INVX2_14 ( .A(A[4]), .Y(_79_) );
NOR2X1 NOR2X1_117 ( .A(B[0]), .B(_79_), .Y(_80_) );
NOR2X1 NOR2X1_118 ( .A(_25_), .B(_80_), .Y(_81_) );
NAND3X1 NAND3X1_97 ( .A(_679_), .B(_81_), .C(_28_), .Y(_82_) );
OAI21X1 OAI21X1_184 ( .A(_32_), .B(_56_), .C(_79_), .Y(_83_) );
NAND3X1 NAND3X1_98 ( .A(_387__bF_buf2), .B(_82_), .C(_83_), .Y(_84_) );
NOR2X1 NOR2X1_119 ( .A(A[3]), .B(_299__bF_buf2), .Y(_85_) );
INVX2 INVX2_15 ( .A(_85_), .Y(_86_) );
OAI21X1 OAI21X1_185 ( .A(A[4]), .B(_45_), .C(_82_), .Y(_87_) );
NAND2X1 NAND2X1_115 ( .A(B_1_bF_buf3_), .B(_87_), .Y(_88_) );
NAND3X1 NAND3X1_99 ( .A(_84_), .B(_86_), .C(_88_), .Y(_89_) );
NAND3X1 NAND3X1_100 ( .A(_78_), .B(_84_), .C(_89_), .Y(_90_) );
NAND3X1 NAND3X1_101 ( .A(_69_), .B(_77_), .C(_90_), .Y(_91_) );
AOI21X1 AOI21X1_71 ( .A(_91_), .B(_60_), .C(_365_), .Y(_92_) );
OAI21X1 OAI21X1_186 ( .A(_84_), .B(_76_), .C(_78_), .Y(_93_) );
AOI21X1 AOI21X1_72 ( .A(_93_), .B(_69_), .C(_59_), .Y(_94_) );
XOR2X1 XOR2X1_32 ( .A(_87_), .B(B_1_bF_buf2_), .Y(_95_) );
INVX1 INVX1_109 ( .A(_74_), .Y(_96_) );
OAI21X1 OAI21X1_187 ( .A(_32_), .B(_56_), .C(_96_), .Y(_97_) );
NAND3X1 NAND3X1_102 ( .A(_70_), .B(_71_), .C(_45_), .Y(_98_) );
NAND3X1 NAND3X1_103 ( .A(_486__bF_buf3), .B(_97_), .C(_98_), .Y(_99_) );
NAND3X1 NAND3X1_104 ( .A(B_2_bF_buf3_), .B(_73_), .C(_75_), .Y(_100_) );
NAND2X1 NAND2X1_116 ( .A(_100_), .B(_99_), .Y(_101_) );
NAND3X1 NAND3X1_105 ( .A(_101_), .B(_95_), .C(_69_), .Y(_102_) );
OAI21X1 OAI21X1_188 ( .A(_85_), .B(_102_), .C(_94_), .Y(_103_) );
INVX2 INVX2_16 ( .A(A[3]), .Y(_104_) );
NAND2X1 NAND2X1_117 ( .A(_299__bF_buf1), .B(_104_), .Y(_105_) );
NOR2X1 NOR2X1_120 ( .A(_299__bF_buf0), .B(_104_), .Y(_106_) );
INVX1 INVX1_110 ( .A(_106_), .Y(_107_) );
endmodule
